----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:31:14 01/29/2014 
-- Design Name: 
-- Module Name:    atlys_lab_video - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity atlys_lab_video is
    port ( 
             clk   : in  std_logic; -- 100 MHz
             reset : in  std_logic;
				 SW6   : in  std_logic;
				 up    : in  std_logic;
             down  : in  std_logic;
             tmds  : out std_logic_vector(3 downto 0);
             tmdsb : out std_logic_vector(3 downto 0)
         );
end atlys_lab_video;

-- TODO: Include requied libraries and packages
--       Don't forget about `unisim` and its `vcomponents` package.
-- TODO: Entity declaration (as shown on previous page)

architecture bentley of atlys_lab_video is
    -- TODO: Signals, as needed
	 signal serialize_clk, serialize_clk_n : std_logic;
	 
	 signal pixel_clk, h_sync, v_sync, blank, v_comp : std_logic;
	 
	 signal red_s, green_s, blue_s, clock_s : std_logic;
	 
	 signal red, green, blue : std_logic_vector(7 downto 0);
	 
	 signal row_sig, col_sig : unsigned(10 downto 0);
	 
	 signal ball_x, ball_y, paddle_y : unsigned(10 downto 0);
begin

    -- Clock divider - creates pixel clock from 100MHz clock
    inst_DCM_pixel: DCM
    generic map(
                   CLKFX_MULTIPLY => 2,
                   CLKFX_DIVIDE   => 8,
                   CLK_FEEDBACK   => "1X"
               )
    port map(
                clkin => clk,
                rst   => reset,
                clkfx => pixel_clk
             );

    -- Clock divider - creates HDMI serial output clock
    inst_DCM_serialize: DCM
    generic map(
                   CLKFX_MULTIPLY => 10, -- 5x speed of pixel clock
                   CLKFX_DIVIDE   => 8,
                   CLK_FEEDBACK   => "1X"
               )
    port map(
                clkin => clk,
                rst   => reset,
                clkfx => serialize_clk,
                clkfx180 => serialize_clk_n
            );

	 vga_inst: entity work.vga_sync(moore)
			port map(
				clk  => pixel_clk,
				reset => reset,
				h_sync => h_sync,
				v_sync => v_sync,
				v_completed => v_comp,
				blank => blank,
				row => row_sig,
				column => col_sig
		   );
	 
    pong_control_inst : entity work.pong_control(moore)
			port map( 
				clk => pixel_clk,
				reset => reset,
				up => up,
				down => down,
				v_completed => v_comp,
				ball_x => ball_x,
				ball_y => ball_y,
				paddle_y => paddle_y
			);
	 
	 pixel_inst: entity work.pixel_gen(sel_arch)
			port map(
				row => row_sig, 
				column => col_sig, 
				blank => blank,
				switch_6 => SW6,
				ball_x => ball_x,
				ball_y =>  ball_y,
				paddle_y => paddle_y,
				r => red, 
				g => green, 
				b => blue
			);

    -- Convert VGA signals to HDMI (actually, DVID ... but close enough)
    inst_dvid: entity work.dvid
    port map(
                clk       => serialize_clk,
                clk_n     => serialize_clk_n, 
                clk_pixel => pixel_clk,
                red_p     => red,
                green_p   => green,
                blue_p    => blue,
                blank     => blank,
                hsync     => h_sync,
                vsync     => v_sync,
                -- outputs to TMDS drivers
                red_s     => red_s,
                green_s   => green_s,
                blue_s    => blue_s,
                clock_s   => clock_s
            );

    -- Output the HDMI data on differential signalling pins
    OBUFDS_blue  : OBUFDS port map
        ( O  => TMDS(0), OB => TMDSB(0), I  => blue_s  );
    OBUFDS_red   : OBUFDS port map
        ( O  => TMDS(1), OB => TMDSB(1), I  => green_s );
    OBUFDS_green : OBUFDS port map
        ( O  => TMDS(2), OB => TMDSB(2), I  => red_s   );
    OBUFDS_clock : OBUFDS port map
        ( O  => TMDS(3), OB => TMDSB(3), I  => clock_s );

end bentley;